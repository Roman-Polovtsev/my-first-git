module verilog_git
(
    input logic a
);
 always_comb
   begin
       a= 1;
   end
endmodule