module submodule
(
    output logic c
);

always_latch
begin
    c= 0;
end

endmodule